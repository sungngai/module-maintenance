library verilog;
use verilog.vl_types.all;
entity pllnrst_vlg_tst is
end pllnrst_vlg_tst;
